library ieee;
use ieee.std_logic_1164.all;

entity LFSR10Test is
end entity LFSR10Test;
 
architecture Behavioural of LFSR10Test is
	constant ClockPeriod : time := 5 ms;
	signal Clock : std_ulogic := '0';
	signal Shift : std_ulogic := '0';
	signal Reset : std_ulogic := '0';
	signal Data : std_ulogic;
begin
	uut : entity work.LFSR10
	port map(
		Clock => Clock,
		Shift => Shift,
		Reset => Reset,
		Data => Data
	);

	process
		procedure Tick is
		begin
			wait for ClockPeriod / 4;
			Clock <= '1';
			wait for ClockPeriod / 2;
			Clock <= '0';
			wait for ClockPeriod / 4;
		end procedure Tick;
	begin
		Tick;
		assert Data = '1';
		Shift <= '1';

		-- This was autogenerated to test that the 1024-bit sequence is
		-- equivalent to a 1024-bit sequence generated by a C program that
		-- ostensibly implemented the same LFSR.
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '0';
		Tick;
		assert Data = '1';
		Tick;
		assert Data = '1';

		wait;
	end process;
end architecture Behavioural;
