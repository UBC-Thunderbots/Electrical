package commands is
	constant COMMAND_READ_DNA : natural := 16#00#;
	constant COMMAND_READ_SWITCHES : natural := 16#01#;
	constant COMMAND_WRITE_LEDS : natural := 16#02#;
	constant COMMAND_GET_CLEAR_IRQS : natural := 16#10#;
	constant COMMAND_MRF_DA_READ_SHORT : natural := 16#20#;
	constant COMMAND_MRF_DA_WRITE_SHORT : natural := 16#21#;
	constant COMMAND_MRF_DA_READ_LONG : natural := 16#22#;
	constant COMMAND_MRF_DA_WRITE_LONG : natural := 16#23#;
	constant COMMAND_MRF_DA_GET_DATA : natural := 16#24#;
	constant COMMAND_MRF_DA_GET_INT : natural := 16#25#;
	constant COMMAND_MRF_DA_SET_AUX : natural := 16#26#;
	constant COMMAND_MRF_OFFLOAD : natural := 16#27#;
	constant COMMAND_MRF_RX_GET_SIZE : natural := 16#28#;
	constant COMMAND_MRF_RX_READ : natural := 16#29#;
	constant COMMAND_MRF_TX_PUSH : natural := 16#2A#;
	constant COMMAND_MRF_TX_GET_STATUS : natural := 16#2B#;
	constant COMMAND_MRF_OFFLOAD_DISABLE : natural := 16#2C#;
	constant COMMAND_MOTORS_SET : natural := 16#30#;
	constant COMMAND_MOTORS_GET_HALL_COUNT : natural := 16#31#;
	constant COMMAND_MOTORS_GET_CLEAR_STUCK_HALLS : natural := 16#32#;
	constant COMMAND_SENSORS_GET_ACCEL : natural := 16#40#;
	constant COMMAND_SENSORS_GET_GYRO : natural := 16#41#;
end package commands;
