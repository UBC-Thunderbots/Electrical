library ieee;
use ieee.std_logic_1164.all;

entity XBeeByteReceiver is
	port(
		Clock1 : in std_ulogic;

		SerialData : in std_ulogic_vector(7 downto 0);
		SerialStrobe : in std_ulogic;

		Data : out std_ulogic_vector(7 downto 0) := X"00";
		Strobe : out std_ulogic := '0';
		SOP : out std_ulogic := '0'
	);
end entity XBeeByteReceiver;

architecture Behavioural of XBeeByteReceiver is
	signal Escaped : boolean := false;
begin
	Data <= SerialData xor X"20" when Escaped else SerialData;
	Strobe <= '1' when SerialStrobe = '1' and SerialData /= X"7D" and SerialData /= X"7E" else '0';
	SOP <= '1' when SerialStrobe = '1' and SerialData = X"7E" else '0';

	process(Clock1)
	begin
		if rising_edge(Clock1) then
			if SerialStrobe = '1' then
				if SerialData = X"7D" then
					Escaped <= true;
				else
					Escaped <= false;
				end if;
			end if;
		end if;
	end process;
end architecture Behavioural;
