library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Types.all;

--
-- Implements the control logic.
--
-- This is implemented as a state machine that iterates through a number of states.
-- Each state selects 3 variables, associates them with 3 coefficients, multiplies
-- the coefficients by the variables, adds the products, and stores the result into
-- a variable. At the rising edge of the 100MHz clock, the following happens:
--
-- (1) The computed output of the previous state is latched onto the appropriate variable.
-- (2) The state variable takes on the appropriate value.
-- (2a) This causes the variables to be multiplied are muxed into the multipliers.
-- (3) The ROMs present the coefficients to the multipliers.
-- (4) The address inputs to the ROMs take on the address for the next clock edge.
--
-- Between that rising edge and the next edge, the MAdd computes the output for the inputs.
--
entity Controller is
	port(
		Clock1 : in std_ulogic;
		Clock100 : in std_ulogic;

		ControlledDriveFlag : in std_ulogic;
		VelocitiesFlag : in std_ulogic;

		Drive1 : in signed(15 downto 0);
		Drive2 : in signed(15 downto 0);
		Drive3 : in signed(15 downto 0);
		Drive4 : in signed(15 downto 0);

		Encoder1 : in signed(17 downto 0);
		Encoder2 : in signed(17 downto 0);
		Encoder3 : in signed(17 downto 0);
		Encoder4 : in signed(17 downto 0);

		Motor1 : out signed(10 downto 0);
		Motor2 : out signed(10 downto 0);
		Motor3 : out signed(10 downto 0);
		Motor4 : out signed(10 downto 0)
	);
end entity Controller;

architecture Behavioural of Controller is
	signal ROMAddress : natural range 0 to 7;
	signal Coeff1Raw : std_ulogic_vector(17 downto 0);
	signal Coeff2Raw : std_ulogic_vector(17 downto 0);
	signal Coeff3Raw : std_ulogic_vector(17 downto 0);

	signal Coeff1 : signed(17 downto 0);
	signal Coeff2 : signed(17 downto 0);
	signal Coeff3 : signed(17 downto 0);
	signal Var1 : signed(17 downto 0);
	signal Var2 : signed(17 downto 0);
	signal Var3 : signed(17 downto 0);
	signal Prod : signed(35 downto 0);

	signal V2MOut1 : signed(35 downto 0);
	signal V2MOut2 : signed(35 downto 0);
	signal V2MOut3 : signed(35 downto 0);
	signal V2MOut4 : signed(35 downto 0);

	signal Setpoint1 : signed(17 downto 0);
	signal Setpoint2 : signed(17 downto 0);
	signal Setpoint3 : signed(17 downto 0);
	signal Setpoint4 : signed(17 downto 0);

	signal Error1 : signed(17 downto 0);
	signal Error2 : signed(17 downto 0);
	signal Error3 : signed(17 downto 0);
	signal Error4 : signed(17 downto 0);

	type StateType is (V2M1, V2M2, V2M3, V2M4, PID1, PID2, PID3, PID4);
	pure function NextState(State : StateType) return StateType is
	begin
		if State = V2M1 then
			return V2M2;
		elsif State = V2M2 then
			return V2M3;
		elsif State = V2M3 then
			return V2M4;
		elsif State = V2M4 then
			return PID1;
		elsif State = PID1 then
			return PID2;
		elsif State = PID2 then
			return PID3;
		elsif State = PID3 then
			return PID4;
		else
			return V2M1;
		end if;
	end function NextState;

	-- This is the state that's currently displayed in the output latch of the multiplier.
	-- On the next rising edge, it will be captured into the appropriate destination variable.
	signal LatchOutputState : StateType := V2M1;

	-- This is the state that's currently latched in the input latches of the multipliers and
	-- being multiplied.
	signal LatchInputState : StateType;

	-- This is the state whose variables are being muxed into the inputs for latching at the next
	-- clock cycle.
	signal MuxInputState : StateType;

	-- This is the state whose coefficients are currently addressed in the ROMs.
	signal ROMAddressState : StateType;
begin
	-- If some state is latched in the output of the multipliers, then the next state must be
	-- latched in the input of the multipliers and be being multiplied right now.
	LatchInputState <= NextState(LatchOutputState);

	-- If some state is latched in the input of the multipliers, then the next state's variables
	-- should be being routed into the latches for capture on the next clock edge.
	MuxInputState <= NextState(LatchInputState);

	-- If some state's variables and coefficients are being routed into the multipliers, then the
	-- coefficients for that state are in the output latches of the ROMs. The ROMs' address inputs
	-- should be seeing the address for the next state, so that on the next rising edge, the data
	-- at that address will appear on the ROM outputs.
	ROMAddressState <= NextState(MuxInputState);

	MAddInstance : entity work.MAdd(Behavioural)
	port map(
		Clock => Clock100,
		A => Coeff1,
		B => Coeff2,
		C => Coeff3,
		X => Var1,
		Y => Var2,
		Z => Var3,
		Prod => Prod
	);
	Coeffs1 : entity work.ROM(Behavioural)
	generic map(
		InitData =>
		(
			-- First **column** of V2M matrix.
			std_ulogic_vector(to_signed(1, 18)),
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(0, 18)),
			-- Proportional coefficients for motors 1, 2, 3, 4.
			std_ulogic_vector(to_signed(1, 18)),
			std_ulogic_vector(to_signed(1, 18)),
			std_ulogic_vector(to_signed(1, 18)),
			std_ulogic_vector(to_signed(1, 18))
		)
	)
	port map(
		Clock => Clock100,
		Address => ROMAddress,
		Data => Coeff1Raw
	);
	Coeffs2 : entity work.ROM(Behavioural)
	generic map(
		InitData =>
		(
			-- Second **column** of V2M matrix.
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(1, 18)),
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(0, 18)),
			-- Integral coefficients for motors 1, 2, 3, 4.
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(0, 18))
		)
	)
	port map(
		Clock => Clock100,
		Address => ROMAddress,
		Data => Coeff2Raw
	);
	Coeffs3 : entity work.ROM(Behavioural)
	generic map(
		InitData =>
		(
			-- Third **column** of V2M matrix.
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(1, 18)),
			std_ulogic_vector(to_signed(0, 18)),
			-- Derivative coefficients for motors 1, 2, 3, 4.
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(0, 18)),
			std_ulogic_vector(to_signed(0, 18))
		)
	)
	port map(
		Clock => Clock100,
		Address => ROMAddress,
		Data => Coeff3Raw
	);
	Coeff1 <= signed(Coeff1Raw);
	Coeff2 <= signed(Coeff2Raw);
	Coeff3 <= signed(Coeff3Raw);

	-- The PID loops take their inputs either from the outputs of the matrix or
	-- from the drive values directly, depending on the flags.
	process(ControlledDriveFlag, VelocitiesFlag, Drive1, Drive2, Drive3, Drive4, V2MOut1, V2MOut2, V2MOut3, V2MOut4)
	begin
		if ControlledDriveFlag = '1' then
			Setpoint1 <= resize(Drive1, Setpoint1'length);
			Setpoint2 <= resize(Drive2, Setpoint2'length);
			Setpoint3 <= resize(Drive3, Setpoint3'length);
			Setpoint4 <= resize(Drive4, Setpoint4'length);
		elsif VelocitiesFlag = '1' then
			Setpoint1 <= V2MOut1(17 downto 0);
			Setpoint2 <= V2MOut2(17 downto 0);
			Setpoint3 <= V2MOut3(17 downto 0);
			Setpoint4 <= V2MOut4(17 downto 0);
		else
			Setpoint1 <= to_signed(0, 18);
			Setpoint2 <= to_signed(0, 18);
			Setpoint3 <= to_signed(0, 18);
			Setpoint4 <= to_signed(0, 18);
		end if;
	end process;

	-- PID uses errors, which are differences between setpoints and encoder-provided plant values.
	Error1 <= Setpoint1 - Encoder1;
	Error2 <= Setpoint2 - Encoder2;
	Error3 <= Setpoint3 - Encoder3;
	Error4 <= Setpoint4 - Encoder4;

	-- Depending on the state, we must select the proper address for the ROMs.
	ROMAddress <=
		     0 when ROMAddressState = V2M1
		else 1 when ROMAddressState = V2M2
		else 2 when ROMAddressState = V2M3
		else 3 when ROMAddressState = V2M4
		else 4 when ROMAddressState = PID1
		else 5 when ROMAddressState = PID2
		else 6 when ROMAddressState = PID3
		else 7 when ROMAddressState = PID4;

	-- Depending on the state, we must select the proper inputs to the MAdd.
	process(MuxInputState, Drive1, Drive2, Drive3, Error1, Error2, Error3, Error4)
	begin
		if MuxInputState = V2M1 then
			Var1 <= resize(Drive1, Var1'length);
			Var2 <= resize(Drive2, Var2'length);
			Var3 <= resize(Drive3, Var3'length);
		elsif MuxInputState = V2M2 then
			Var1 <= resize(Drive1, Var1'length);
			Var2 <= resize(Drive2, Var2'length);
			Var3 <= resize(Drive3, Var3'length);
		elsif MuxInputState = V2M3 then
			Var1 <= resize(Drive1, Var1'length);
			Var2 <= resize(Drive2, Var2'length);
			Var3 <= resize(Drive3, Var3'length);
		elsif MuxInputState = V2M4 then
			Var1 <= resize(Drive1, Var1'length);
			Var2 <= resize(Drive2, Var2'length);
			Var3 <= resize(Drive3, Var3'length);
		elsif MuxInputState = PID1 then
			Var1 <= Error1;
			Var2 <= to_signed(0, 18);
			Var3 <= to_signed(0, 18);
		elsif MuxInputState = PID2 then
			Var1 <= Error2;
			Var2 <= to_signed(0, 18);
			Var3 <= to_signed(0, 18);
		elsif MuxInputState = PID3 then
			Var1 <= Error3;
			Var2 <= to_signed(0, 18);
			Var3 <= to_signed(0, 18);
		elsif MuxInputState = PID4 then
			Var1 <= Error4;
			Var2 <= to_signed(0, 18);
			Var3 <= to_signed(0, 18);
		end if;
	end process;

	-- On a clock edge, capture the computed output and advance the state variable.
	process(Clock100)
	begin
		if rising_edge(Clock100) then
			if LatchOutputState = V2M1 then
				V2MOut1 <= Prod;
			elsif LatchOutputState = V2M2 then
				V2MOut2 <= Prod;
			elsif LatchOutputState = V2M3 then
				V2MOut3 <= Prod;
			elsif LatchOutputState = V2M4 then
				V2MOut4 <= Prod;
			elsif LatchOutputState = PID1 then
				Motor1 <= Prod(10 downto 0);
			elsif LatchOutputState = PID2 then
				Motor2 <= Prod(10 downto 0);
			elsif LatchOutputState = PID3 then
				Motor3 <= Prod(10 downto 0);
			elsif LatchOutputState = PID4 then
				Motor4 <= Prod(10 downto 0);
			end if;
			LatchOutputState <= NextState(LatchOutputState);
		end if;
	end process;
end architecture Behavioural;
