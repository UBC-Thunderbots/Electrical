library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Types is
	type ROMDataType is array(natural range <>) of std_ulogic_vector(17 downto 0);
end package Types;
